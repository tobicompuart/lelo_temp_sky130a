*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/LELO_TEMP_lpe.spi
#else
.include ../../../work/xsch/LELO_TEMP.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3
*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

.param fLfClk = 32678
.param PERIOD_CLK = 1/fLfClk
.param PW_CLK = PERIOD_CLK/2
*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
VLFCLK lfClk 0 dc 0 pulse (0 {AVDD} 0 {TRF} {TRF} {PW_CLK} {PERIOD_CLK})
VSTART  start  VSS  pwl 0 0 {t_start} 0 {{t_start} + 10p} {AVDD}

Vrst_n rst_n 0 dc {AVDD}

R3 PWRUP_1V8 VDD_1V8 10k
R1 pwrupOsc PWRUP_1V8 1
R2 clk OSC_TEMP_1V8 1

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi
*.include ../svinst_tc.spi
.include ../svinst_tfsm.spi
*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
*.save all
.save v(vdd_1v8) v(vss) v(pwrup_1v8) v(osc_temp_1v8)
.save v(xdut.LPI) v(xdut.CMPO) v(xdut.clk)
.save i(vdd) v(xdut.ibp_1u<0>) v(xdut.vc) v(xdut.rst)
.save v(xdut.x1_ibp.vr1) v(xdut.x1_ibp.vd2)
.save v(lfClk) v(rst_n) v(start)

#ifdef Debug
.option savecurrents
.save all
#endif
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

*- Override the default digital output bridge.
pre_set auto_bridge_d_out =
     + ( ".model auto_dac dac_bridge(out_low = 0.0 out_high = 1.8)"
     +   "auto_bridge%d [ %s ] [ %s ] auto_dac" )

optran 0 0 0 1n 1u 0

tran 1n {t_stop}

write

quit


.endc

.end
