*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/LELO_TEMP_lpe.spi
#else
.include ../../../work/xsch/LELO_TEMP.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-4
.option TEMP=-40
.option TEMP=125
*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
VPWR  PWRUP_1V8  VSS  pwl 0 0 1u 0 {1u + 10p} {AVDD}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
*.save all
.save v(vdd_1v8) v(vss) v(pwrup_1v8) v(osc_temp_1v8)
.save v(xdut.LPI) v(xdut.CMPO) v(xdut.clk)
.save i(vdd)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0

#ifdef Nosweep
tran 0.1n {t_stop}
write {cicname}.raw
#else
set fend = .raw
foreach vtemp {temperatures}
  option temp=$vtemp
  tran 0.1n {t_stop}
  write {cicname}_$vtemp$fend
end

#endif

quit


.endc

.end
